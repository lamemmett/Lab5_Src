module userIO(clock, reset, dataIn, enable, requestComplete, dataOut);

endmodule 

module userIO_testbench();
	
endmodule 